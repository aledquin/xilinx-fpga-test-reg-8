/*  contador4.v
    m�dulo cont4
    Contador de 4 bits sin carga paralela
	Tiene salida Enext = 1 si Cuenta=4'hF.
*/

module cont4(	output reg [3:0] Cuenta,	// Valor del contador s�ncrono
				output reg Enext,			// Cuenta == 4'hF => Enext = 1
                input nR,					// Reset negativo as�ncrono
                input E,					// Enabled E=0 deshabilitado, E=1 habilitado
                input CK					// Clock posedge
);

parameter STD_DELAY = 2;
reg [3:0] CuentaR;

// C�lculo as�ncrono del estado siguiente.
// Lista de sensibilidad depende de estado
// actual y variables de control.
// No depende del reloj.
  always @ (Cuenta, E) begin
  if(E==1) begin
	CuentaR = Cuenta + 1;
	Enext = (Cuenta == 4'hF) ? 1: 0;
	end
  end // always as�ncrono
  
// Actualizaci�n s�ncrona del estado
// Reset debe estar inactivo.
// Enable debe estar activo.
// Se actualiza con posedge.
  always @ ( negedge nR, posedge CK )
  begin
    if(nR == 0) begin						// Aqu� se hace reset
		#(STD_DELAY) Cuenta = 0;
		CuentaR = 0;
		Enext = 0;
	end
    else if( E == 1) begin					// Tiene que estar habilitado para contar
      #(STD_DELAY) Cuenta = CuentaR;		// Actualiza estado
	end
end // always s�ncrono

// En este caso la salida de la m�quina es el estado actual.
// No es necesario actualizar la salida.

endmodule
